module decoder_bit (
    input enable,
    output Y
);
    assign Y = enable;
endmodule
